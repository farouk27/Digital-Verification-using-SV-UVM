module SPI_MONITOR(spi_wrapper_interface.MONITOR w_if);

initial begin 
	$monitor("display all the signals");
end

endmodule 


