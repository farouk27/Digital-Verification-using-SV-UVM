module RAM_MONITOR(RAM_if.MONITOR r_if);

initial begin 
	$monitor("display all the signals");
end
endmodule 

