package shared_pkg;
bit	test_finished;

integer	error_count	= 0;
integer	correct_count	= 0;
endpackage
